module str_03;
  string A=("DESIGN_ENGINEER");
  initial begin
    $display("your's output str_03 on A=%s",A.tolower);
  end
endmodule

result
KERNEL: your's output str_03 on A=design_engineer
