class array;
  rand longint print[1:0][2:0][3:0];
endclass


module tb;
  array a1;
  initial begin
    a1=new();
    for(int i=0;i<=8;i++)begin
      $display("value of 2DIMENTIONAL PACKED ARRAY=[%0p]INDEX=[%0d]",a1.print,i);
      a1.randomize();
    end
    
  end
endmodule


Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Sep 22 09:53 2025
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}, '{'{0, 0, 0, 0}, '{0, 0, 0, 0}, '{0, 0, 0, 0}}} ]INDEX=[0]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{-6842783759417550919, -5726203078114608985, -3506964679157472868, 7624370432706573369}, '{-217367992281279212, -8665355824280435118, -220038429141070629, -30574626034906519}, '{-6702453455987789159, -7745529651938689768, 9199369429609243629, 6941540621650691320}}, '{'{-8482030383469778188, 1343846956935585923, -8230982918858637498, -853518915812920572}, '{-2053584789603162183, 459968098334072856, -5775316183779965922, -2144138228187202489}, '{3266198812699807420, -4221798284927248979, 8571759553769747650, -1002023458822650226}}} ]INDEX=[1]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{5297240865832474715, 8512271973111419274, 4789870128884935381, 214265737261407082}, '{7431014241800143053, -1774225655010308327, 4699146087223598463, 3959689045809846111}, '{8553638632450006887, 7519222227742765980, 4966288974572368959, 889881922114504512}}, '{'{4115554587165018363, 6966853592658604903, 1566400497065484844, -6019401131944120654}, '{698448649948967712, -7823242434269072655, -8316465029302650513, -388000363206296604}, '{-8571702172288861854, 408362218456221536, -5133450303789835654, -5364914133146902116}}} ]INDEX=[2]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{-1192650888000470214, -5507249447573693133, 4237039528035788570, 6884408146246385465}, '{7585255089313458516, 3883027210324771201, -8423594568160284177, 2903854434591552032}, '{-1123399577022233167, 8755954158851992513, 7380702733103247375, 7596478095052978741}}, '{'{-5467299252135809038, -894407498621524129, -6601777247260041079, 7653237004266199775}, '{8042941777719416302, -1706490477296601908, -6600395757235063027, 564192086599632073}, '{-3614144819334575685, 852228003441528463, 5295516546194740551, -8986385753419600700}}} ]INDEX=[3]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{-6167207643120870393, -5848277173853885095, -7024125897722267056, 5047328158663011868}, '{6310671979593353694, -111855646927377385, -207682369991487730, 2069631266512661582}, '{-8944389433963439696, 4283819347868299911, -8031807529340898860, 5642412399645858856}}, '{'{-8527706724674577189, 702763971065346006, -865080045963947127, -8486456397039718938}, '{899716880255270117, 3732833887141525373, -3874955940325486622, -5665669694323908918}, '{-5259926823679032622, 1031625552889340084, 6508003801234328279, 8800799832137521422}}} ]INDEX=[4]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{-6239274059912852512, -955418512444846748, -9087021327781343367, -3356641520684299794}, '{-8115236163374133064, 4884405496062227487, -5916154001830605483, -4625285281409554520}, '{2467616445879805213, 6605739298012439451, -3251258406812388758, -1473152937576010115}}, '{'{430397137958967746, -8106292499132806133, 5377333165287706398, -6711917400274508885}, '{2949273574334916424, -1454813990736287568, 8962339026737019585, 1490645203238023342}, '{-5223872858965899749, -3874306635808479526, 3807031234628663409, -9156136109924615542}}} ]INDEX=[5]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{644555526888659411, 6851366128790476848, 3081647741077274353, 8159223490315394481}, '{1297823778633941377, 7388917145622766583, -7467126157872850629, -5400522629545780422}, '{-7954744276241576027, -478045452360443520, 8732979814354254403, 3360062024825508340}}, '{'{-1679270770998194113, 8492277185170019230, 253164961118349248, -4427106590660833780}, '{6202603819904668406, -3402620327336226547, -1088071231418389251, 3272028205600873267}, '{-4974205411279297174, 7423195890962151667, 6033357598910258975, 7428177996216225144}}} ]INDEX=[6]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{7799135164486699050, -3766579962276177427, 4652186175042698409, -3700062954029838952}, '{-4475103976859202080, -2861400230671707832, 6722929367355544283, 1906920868890047524}, '{7841285894274416134, 131574119626302792, -6499875120456330950, -5650337743769800439}}, '{'{6395749372169759816, -7346168777938560107, -1979502270115553372, 5619826101446913273}, '{4517803518701764769, -7958598308726822337, 8787510793588549541, -6875750644904069235}, '{-7738439543282937521, -3298556091003576104, -2518874332471807834, 8836478662730116294}}} ]INDEX=[7]
value of 2DIMENTIONAL PACKED ARRAY=['{'{'{-1523412329394655245, 3939016738372780849, -4843176191067728190, 694136920240348026}, '{-9135697072988980067, -7446663679560240687, -967563463545928323, 346714462365738877}, '{997760950723981510, -1242602297636080249, 3439052709870216928, 592011251700678538}}, '{'{-5573381839688542737, -8811730707531722139, -1862277788682832752, -1149350093581436056}, '{2799105507906828640, -6950980431688850550, -1364437382461335917, -7849970821017222694}, '{-8245963424882333816, 2593836489773689784, -3924395431954962839, -175463309153889817}}} ]INDEX=[8]
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.360 seconds;       Data structure size:   0.0Mb
Mon Sep 22 09:53:36 2025
