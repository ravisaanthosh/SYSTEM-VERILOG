module repeat_loop_95;
  initial begin
    repeat(5)begin
      $display("Trust your own process it's make a time but trust it.............");
      $display("design and verification engineer..");
    end
  end
endmodule

Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug  5 09:06 2025
Trust your own process it's make a time but trust it.............
design and verification engineer.............
Trust your own process it's make a time but trust it.............
design and verification engineer.............
Trust your own process it's make a time but trust it.............
design and verification engineer.............
Trust your own process it's make a time but trust it.............
design and verification engineer.............
Trust your own process it's make a time but trust it.............
design and verification engineer.............
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.460 seconds;       Data structure size:   0.0Mb
Tue Aug  5 09:06:29 2025
Done
      
