module str_07;
  string A="DESIGN 1245";
  initial begin
    $display("your's expected output for str_07 is A=%s",A.itoa());
  end
endmodule

result tool error
work = /home/runner/work/work.lib
ERROR VCP7292 "String method itoa is not a function." 

expected output..!
DESIGN
