module reg_27;
   reg reg_27;
  initial begin
    $display("reg_27=%b",reg_27);
    reg_27 =1'b0;
    $display("reg_27=%b",reg_27);
  end
endmodule
