module byte_28;
   byte byte_28;
  initial begin
    $display("byte_28=%b",byte_28);
    byte_28 =8'b11111111;
    $display("byte_28=%b",byte_28);
  end
endmodule
