module r_26;
   real r_26;
  initial begin
    $display("r__26=%b",r_26);
    r_26 =64'b10101010101011111010;
    $display("r_26=%b",r_26);
  end
endmodule
