  integer int_24;
  initial begin
    $display("int_24=%b",int_24);
    int_24 =4'b1010;
    $display("int_24=%b",int_24);
  end
endmodule
