module str_1;
  string A="DESIGN ENGINEER";
  initial begin
    $display("output A=%d",A.len);
  end
endmodule


expected output_str_1
KERNEL: output A= 15
