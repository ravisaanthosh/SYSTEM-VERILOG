module loop_while_90;
  integer i;
  initial begin
    i=0;
    while(i<=6)begin
      $display("your's while_loops_output is=%0d",i);
    i++;
  end
  end
endmodule

your's while_loops_output is=0
your's while_loops_output is=1
your's while_loops_output is=2
your's while_loops_output is=3
your's while_loops_output is=4
your's while_loops_output is=5
your's while_loops_output is=6
           V C S   S i m u l a t i o n   R e p o r t 
Time: 0 ns
CPU Time:      0.490 seconds;       Data structure size:   0.0Mb
Tue Aug  5 02:30:10 2025
