module long_int31;
   shortint long_int_31;
  initial begin
    $display("long_int_31=%b",long_int_31);
    long_int_31 =64'b11111111;
    $display("long_int_31=%b",long_int_31);
  end
endmodule
