module bit_29;
   bit bit_29;
  initial begin
    $display("bit_29=%b",bit_29);
    bit_29 =8'b11111111;
    $display("bit_29=%b",bit_29);
  end
endmodule
