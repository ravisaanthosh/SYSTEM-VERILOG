module i_23;
  integer int_23;
  initial begin
    $display("int_23=%b",int_23);
    int_23=5'b10101;
     $display("int_23=%b",int_23);
  end
endmodule
