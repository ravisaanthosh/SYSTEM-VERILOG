module t_25;
   time t_25;
  initial begin
    $display("int_25=%b",t_25);
    t_25 =4'b1010;
    $display("int_25=%b",t_25);
  end
endmodule
