module for_loop_93;
  shortint loop;
  initial begin
    for(loop=0; loop<=56; loop=loop+2)
      $display("you's for_loop output is =[%0d]",loop);
  end
endmodule

Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Aug  5 08:39 2025
you's for_loop output is =[0]
you's for_loop output is =[2]
you's for_loop output is =[4]
you's for_loop output is =[6]
you's for_loop output is =[8]
you's for_loop output is =[10]
you's for_loop output is =[12]
you's for_loop output is =[14]
you's for_loop output is =[16]
you's for_loop output is =[18]
you's for_loop output is =[20]
you's for_loop output is =[22]
you's for_loop output is =[24]
you's for_loop output is =[26]
you's for_loop output is =[28]
you's for_loop output is =[30]
you's for_loop output is =[32]
you's for_loop output is =[34]
you's for_loop output is =[36]
you's for_loop output is =[38]
you's for_loop output is =[40]
you's for_loop output is =[42]
you's for_loop output is =[44]
you's for_loop output is =[46]
you's for_loop output is =[48]
you's for_loop output is =[50]
you's for_loop output is =[52]
you's for_loop output is =[54]
you's for_loop output is =[56]
